﻿<?xml version="1.0"?>
<ArrayOfQuestion xmlns:xsi="http://www.w3.org/2001/XMLSchema-instance" xmlns:xsd="http://www.w3.org/2001/XMLSchema">
  <Question>
    <text>В Древнем Риме альбомом называли доску, покрытую белым гипсом.</text>
    <trueFalse>true</trueFalse>
  </Question>
  <Question>
    <text>На луну воют только волки-одиночки.</text>
    <trueFalse>false</trueFalse>
  </Question>
  <Question>
    <text>Бамбук самая высокая трава в мире.</text>
    <trueFalse>true</trueFalse>
  </Question>
  <Question>
    <text>Авторучка была изобретена ещё в Древнем Египте?</text>
    <trueFalse>true</trueFalse>
  </Question>
  <Question>
    <text>Совы не могут вращать глазами?</text>
    <trueFalse>true</trueFalse>
  </Question>
  <Question>
    <text>Дети могут слышать более высокие звуки, чем взрослые?</text>
    <trueFalse>true</trueFalse>
  </Question>
  <Question>
    <text>Лось является разновидностью оленя?</text>
    <trueFalse>true</trueFalse>
  </Question>
  <Question>
    <text>Мойву эскимосы сушат и едят вместо хлеба?</text>
    <trueFalse>true</trueFalse>
  </Question>
  <Question>
    <text>Радугу можно увидеть и в полночь?</text>
    <trueFalse>true</trueFalse>
  </Question>
  <Question>
    <text>Утром вы выше ростом, чем вечером?</text>
    <trueFalse>true</trueFalse>
  </Question>
</ArrayOfQuestion>